`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.06.2024 13:22:15
// Design Name: 
// Module Name: Stage2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module Stage2(
    input Enable,
    input [7:0] a0,a1,a2,a3,b0,b1,b2,b3,c0,c1,c2,c3,d0,d1,d2,d3,
    input k0,k1,
    output reg [7:0] w0,w1,w2,w3,x0,x1,x2,x3,y0,y1,y2,y3,z0,z1,z2,z3
    );

always @ (*) begin
if(Enable)begin
    w0 = 8'b0; w1 = 8'b0; w2 = 8'b0; w3 = 8'b0;
    x0 = 8'b0; x1 = 8'b0; x2 = 8'b0; x3 = 8'b0;
    y0 = 8'b0; y1 = 8'b0; y2 = 8'b0; y3 = 8'b0;
    z0 = 8'b0; z1 = 8'b0; z2 = 8'b0; z3 = 8'b0;
    if(~k0&~k1) begin//67452301
        w0 = {a0[6], a0[7], a0[4], a0[5], a0[2], a0[3], a0[0], a0[1]};
        w1 = {a1[6], a1[7], a1[4], a1[5], a1[2], a1[3], a1[0], a1[1]};
        w2 = {a2[6], a2[7], a2[4], a2[5], a2[2], a2[3], a2[0], a2[1]};
        w3 = {a3[6], a3[7], a3[4], a3[5], a3[2], a3[3], a3[0], a3[1]};
        x0 = {b0[6], b0[7], b0[4], b0[5], b0[2], b0[3], b0[0], b0[1]};
        x1 = {b1[6], b1[7], b1[4], b1[5], b1[2], b1[3], b1[0], b1[1]};
        x2 = {b2[6], b2[7], b2[4], b2[5], b2[2], b2[3], b2[0], b2[1]};
        x3 = {b3[6], b3[7], b3[4], b3[5], b3[2], b3[3], b3[0], b3[1]};
        y0 = {c0[6], c0[7], c0[4], c0[5], c0[2], c0[3], c0[0], c0[1]};
        y1 = {c1[6], c1[7], c1[4], c1[5], c1[2], c1[3], c1[0], c1[1]};
        y2 = {c2[6], c2[7], c2[4], c2[5], c2[2], c2[3], c2[0], c2[1]};
        y3 = {c3[6], c3[7], c3[4], c3[5], c3[2], c3[3], c3[0], c3[1]};
        z0 = {d0[6], d0[7], d0[4], d0[5], d0[2], d0[3], d0[0], d0[1]};
        z1 = {d1[6], d1[7], d1[4], d1[5], d1[2], d1[3], d1[0], d1[1]};
        z2 = {d2[6], d2[7], d2[4], d2[5], d2[2], d2[3], d2[0], d2[1]};
        z3 = {d3[6], d3[7], d3[4], d3[5], d3[2], d3[3], d3[0], d3[1]};
    end
    
    else if (k0&~k1) begin //32107654
        w0 = {a0[3], a0[2], a0[1], a0[0], a0[7], a0[6], a0[5], a0[4]};
        w1 = {a1[3], a1[2], a1[1], a1[0], a1[7], a1[6], a1[5], a1[4]};
        w2 = {a2[3], a2[2], a2[1], a2[0], a2[7], a2[6], a2[5], a2[4]};
        w3 = {a3[3], a3[2], a3[1], a3[0], a3[7], a3[6], a3[5], a3[4]};
        x0 = {b0[3], b0[2], b0[1], b0[0], b0[7], b0[6], b0[5], b0[4]};
        x1 = {b1[3], b1[2], b1[1], b1[0], b1[7], b1[6], b1[5], b1[4]};
        x2 = {b2[3], b2[2], b2[1], b2[0], b2[7], b2[6], b2[5], b2[4]};
        x3 = {b3[3], b3[2], b3[1], b3[0], b3[7], b3[6], b3[5], b3[4]};
        y0 = {c0[3], c0[2], c0[1], c0[0], c0[7], c0[6], c0[5], c0[4]};
        y1 = {c1[3], c1[2], c1[1], c1[0], c1[7], c1[6], c1[5], c1[4]};
        y2 = {c2[3], c2[2], c2[1], c2[0], c2[7], c2[6], c2[5], c2[4]};
        y3 = {c3[3], c3[2], c3[1], c3[0], c3[7], c3[6], c3[5], c3[4]};
        z0 = {d0[3], d0[2], d0[1], d0[0], d0[7], d0[6], d0[5], d0[4]};
        z1 = {d1[3], d1[2], d1[1], d1[0], d1[7], d1[6], d1[5], d1[4]};
        z2 = {d2[3], d2[2], d2[1], d2[0], d2[7], d2[6], d2[5], d2[4]};
        z3 = {d3[3], d3[2], d3[1], d3[0], d3[7], d3[6], d3[5], d3[4]};
    end
    else if(~k0&k1) begin // left 2
        w0 = {a0[0], a0[1], a0[2], a0[3], a0[4], a0[5], a0[6], a0[7]};
        w1 = {a1[0], a1[1], a1[2], a1[3], a1[4], a1[5], a1[6], a1[7]};
        w2 = {a2[0], a2[1], a2[2], a2[3], a2[4], a2[5], a2[6], a2[7]};
        w3 = {a3[0], a3[1], a3[2], a3[3], a3[4], a3[5], a3[6], a3[7]};
        x0 = {b0[0], b0[1], b0[2], b0[3], b0[4], b0[5], b0[6], b0[7]};
        x1 = {b1[0], b1[1], b1[2], b1[3], b1[4], b1[5], b1[6], b1[7]};
        x2 = {b2[0], b2[1], b2[2], b2[3], b2[4], b2[5], b2[6], b2[7]};
        x3 = {b3[0], b3[1], b3[2], b3[3], b3[4], b3[5], b3[6], b3[7]};
        y0 = {c0[0], c0[1], c0[2], c0[3], c0[4], c0[5], c0[6], c0[7]};
        y1 = {c1[0], c1[1], c1[2], c1[3], c1[4], c1[5], c1[6], c1[7]};
        y2 = {c2[0], c2[1], c2[2], c2[3], c2[4], c2[5], c2[6], c2[7]};
        y3 = {c3[0], c3[1], c3[2], c3[3], c3[4], c3[5], c3[6], c3[7]};
        z0 = {d0[0], d0[1], d0[2], d0[3], d0[4], d0[5], d0[6], d0[7]};
        z1 = {d1[0], d1[1], d1[2], d1[3], d1[4], d1[5], d1[6], d1[7]};
        z2 = {d2[0], d2[1], d2[2], d2[3], d2[4], d2[5], d2[6], d2[7]};
        z3 = {d3[0], d3[1], d3[2], d3[3], d3[4], d3[5], d3[6], d3[7]};
    end
    else if (k0&k1) begin
        w0 = {a0[1], a0[6], a0[3], a0[4], a0[5], a0[2], a0[7], a0[0]};
        w1 = {a1[1], a1[6], a1[3], a1[4], a1[5], a1[2], a1[7], a1[0]};
        w2 = {a2[1], a2[6], a2[3], a2[4], a2[5], a2[2], a2[7], a2[0]};
        w3 = {a3[1], a3[6], a3[3], a3[4], a3[5], a3[2], a3[7], a3[0]};
        x0 = {b0[1], b0[6], b0[3], b0[4], b0[5], b0[2], b0[7], b0[0]};
        x1 = {b1[1], b1[6], b1[3], b1[4], b1[5], b1[2], b1[7], b1[0]};
        x2 = {b2[1], b2[6], b2[3], b2[4], b2[5], b2[2], b2[7], b2[0]};
        x3 = {b3[1], b3[6], b3[3], b3[4], b3[5], b3[2], b3[7], b3[0]};
        y0 = {c0[1], c0[6], c0[3], c0[4], c0[5], c0[2], c0[7], c0[0]};
        y1 = {c1[1], c1[6], c1[3], c1[4], c1[5], c1[2], c1[7], c1[0]};
        y2 = {c2[1], c2[6], c2[3], c2[4], c2[5], c2[2], c2[7], c2[0]};
        y3 = {c3[1], c3[6], c3[3], c3[4], c3[5], c3[2], c3[7], c3[0]};
        z0 = {d0[1], d0[6], d0[3], d0[4], d0[5], d0[2], d0[7], d0[0]};
        z1 = {d1[1], d1[6], d1[3], d1[4], d1[5], d1[2], d1[7], d1[0]};
        z2 = {d2[1], d2[6], d2[3], d2[4], d2[5], d2[2], d2[7], d2[0]};
        z3 = {d3[1], d3[6], d3[3], d3[4], d3[5], d3[2], d3[7], d3[0]};
    end
  end
else begin
    w0 = 8'bZ; w1 = 8'bZ; w2 = 8'bZ; w3 = 8'bZ;
    x0 = 8'bZ; x1 = 8'bZ; x2 = 8'bZ; x3 = 8'bZ;
    y0 = 8'bZ; y1 = 8'bZ; y2 = 8'bZ; y3 = 8'bZ;
    z0 = 8'bZ; z1 = 8'bZ; z2 = 8'bZ; z3 = 8'bZ;
end
end    
endmodule
// k1   k0   y 
// 0    0    67452301
// 0    1    32107654
// 1    0    01234567
// 1    1    16345270
